interface fifo_if(input bit clk);
    parameter FIFO_WIDTH = 16;
    parameter FIFO_DEPTH = 8;
    logic [FIFO_WIDTH-1:0] data_in;
    logic rst_n; 
    logic wr_en;
    logic rd_en;
    logic  [FIFO_WIDTH-1:0] data_out;
    logic  wr_ack;
    logic overflow;
    logic full, empty, almostfull, almostempty, underflow;
    modport dut(
        input data_in, wr_en, rd_en, clk, rst_n,
        output full, empty, almostfull, almostempty, wr_ack, overflow, underflow, data_out
    );
    modport test(
        output data_in, wr_en, rd_en, rst_n,
        input clk,full, empty, almostfull, almostempty, wr_ack, overflow, underflow, data_out
    );
    modport monitor(
        input data_in, wr_en, rd_en, rst_n,clk,full, empty, almostfull, almostempty, wr_ack, overflow, underflow, data_out
    );


endinterface